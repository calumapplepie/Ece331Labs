* Wey Makeup Calum McConnell
* full disclosure: i restarted from the original Lab1 spice deck, since I was on a new machine

.include Problem5.inc

* Setting up the voltage signal source for DC, AC and Transient Analysis
Vsig Vsig 0 DC 5 AC 1 0 PULSE(0,5,5ms,0.001ms,0.001ms,5ms,10ms)
Vsupply Vsupply 0 DC 5
* Syntax:  Vx + - DC (DCVALUE) AC (ACVALUE) (ACPHASE) (Transient Signal)

* Setup Passive Components
R1 Vsupply Va 540;  10K series resistor
XLED Va Vc LED
Mx Vc Vsig 0 0 CMOSN W=41.67u L=1u

* Setup simulation temperature in Celsius
.TEMP 25C

* Setup DC Analysis
*.DC Vsig -5 5 0.1 ; Syntax .DC Source Vstart Vstop Vstep
* Alternatively the statement .DC Vsig 5 -5 -0.1 will go from 5V to -5V in -0.1V steps
* DC Analysis: Spice will vary the DC value of the declared swept source.  All other sources held at their DC values.

* Setup AC Analysis
*.AC DEC 20 100 10K ; Syntax: .AC (LIN/OCT/DEC) Points Fstart Fstop
* You must declare all values.
* AC Analysis: Spice first performs an operating point calculation at the DC declared value of Vsig and Iload
* and then performs an AC analysis using only the AC declared values.  Note this is a frequency domain (jw) and superposition technique,
* the AC analysis results are due only to the AC inputs.
* Note: Typically we will only evaluate 1 AC source at a time.

* Transient Analysis
.TRAN 1ms 30mS 0 0.1ms ; Syntax: .TRAN Printstep StopTime PrintStartTime MaximumStepSize
* You must declare Printstep and simulation stoptime.
* Transient Analysis:  In transient analysis, Spice ignores the AC declaration and only uses the DC declaration
* if no transient declaration exists.  To begin the simulation, Spice performs a bias point calculation time=0.

* Probe Statement - Generates .PRB file for Post Processor, your Spice file should include it
.Probe
*
.End

* Good practice to use a .end card although some spice simulators don't need it.







